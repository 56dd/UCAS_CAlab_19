module div(
    
);

endmodule