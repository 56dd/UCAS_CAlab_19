module mul(
    
);

endmodule